VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO project1
  CLASS BLOCK ;
  FOREIGN project1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 34.500 BY 57.120 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.020 10.640 14.620 46.480 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 10.640 11.320 46.480 ;
    END
  END VPWR
  PIN in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END in1[0]
  PIN in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END in1[1]
  PIN in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END in1[2]
  PIN in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END in1[3]
  PIN in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END in1[4]
  PIN in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END in1[5]
  PIN in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END in1[6]
  PIN in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END in1[7]
  PIN out1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 30.500 51.720 34.500 52.320 ;
    END
  END out1[0]
  PIN out1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 30.500 44.920 34.500 45.520 ;
    END
  END out1[1]
  PIN out1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 30.500 38.120 34.500 38.720 ;
    END
  END out1[2]
  PIN out1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 30.500 31.320 34.500 31.920 ;
    END
  END out1[3]
  PIN out1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 30.500 24.520 34.500 25.120 ;
    END
  END out1[4]
  PIN out1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 30.500 17.720 34.500 18.320 ;
    END
  END out1[5]
  PIN out1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 30.500 10.920 34.500 11.520 ;
    END
  END out1[6]
  PIN out1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 30.500 4.120 34.500 4.720 ;
    END
  END out1[7]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 29.170 46.430 ;
      LAYER li1 ;
        RECT 5.520 10.795 28.980 46.325 ;
      LAYER met1 ;
        RECT 4.210 10.640 28.980 46.480 ;
      LAYER met2 ;
        RECT 4.230 4.235 27.510 52.205 ;
      LAYER met3 ;
        RECT 4.400 51.320 30.100 52.185 ;
        RECT 3.990 45.920 30.500 51.320 ;
        RECT 4.400 44.520 30.100 45.920 ;
        RECT 3.990 39.120 30.500 44.520 ;
        RECT 4.400 37.720 30.100 39.120 ;
        RECT 3.990 32.320 30.500 37.720 ;
        RECT 4.400 30.920 30.100 32.320 ;
        RECT 3.990 25.520 30.500 30.920 ;
        RECT 4.400 24.120 30.100 25.520 ;
        RECT 3.990 18.720 30.500 24.120 ;
        RECT 4.400 17.320 30.100 18.720 ;
        RECT 3.990 11.920 30.500 17.320 ;
        RECT 4.400 10.520 30.100 11.920 ;
        RECT 3.990 5.120 30.500 10.520 ;
        RECT 4.400 4.255 30.100 5.120 ;
      LAYER met4 ;
        RECT 25.135 12.415 25.465 35.185 ;
  END
END project1
END LIBRARY

